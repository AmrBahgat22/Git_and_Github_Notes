library verilog;
use verilog.vl_types.all;
entity Parity_Generator_Tx_tb is
end Parity_Generator_Tx_tb;

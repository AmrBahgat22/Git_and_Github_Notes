library verilog;
use verilog.vl_types.all;
entity PISO_Register_tb is
end PISO_Register_tb;

library verilog;
use verilog.vl_types.all;
entity Baud_Rate_Generator_Tx_tb is
end Baud_Rate_Generator_Tx_tb;

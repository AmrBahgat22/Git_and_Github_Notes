library verilog;
use verilog.vl_types.all;
entity Transmitter_FSM_tb is
end Transmitter_FSM_tb;
